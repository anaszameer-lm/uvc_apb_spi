package apb_package;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "tb_src/apb_transaction.sv"
`include "tb_src/apb_sequence.sv" 
`include "tb_src/apb_sequencer.sv"
`include "tb_src/apb_driver.sv"
`include "tb_src/apb_monitor.sv"
`include "tb_src/apb_agent.sv"
`include "tb_src/apb_scoreboard.sv"    
`include "tb_src/apb_environment.sv"
`include "tb_src/apb_test.sv"    


endpackage : apb_package
